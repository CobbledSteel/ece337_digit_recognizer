
`timescale 1ns / 10ps

module tb_sigmoid_ALU ();

endmodule
