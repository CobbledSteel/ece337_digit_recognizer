// $Id: $
// File name:   stp_shift_reg.sv
// Created:     4/4/2018
// Author:      Chan Weng Yan
// Lab Section: 337-08
// Version:     1.0  Initial Design Entry
// Description: Serial-to-parallel shift register
