// $Id: $
// File name:   tb_digit_recognizer.sv
// Created:     4/21/2018
// Author:      Group
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Top level testbench for digit recognizer
