// $Id: $
// File name:   spi_input.sv
// Created:     4/20/2018
// Author:      Chan Weng Yan
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: SPI input controller file

