// $Id: $
// File name:   tb_digit_recognizer.sv
// Created:     4/21/2018
// Author:      Chan Weng Yan
// Lab Section: 337-08
// Version:     1.0  Initial Design Entry
// Description: Top level testbench for digit recognizer
