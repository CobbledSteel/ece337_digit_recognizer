// $Id: $
// File name:   sigmoid_ALU_signed_adder.sv
// Created:     4/4/2018
// Author:      Vadim Nikiforov
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: signed adder for the sigmoid ALU
