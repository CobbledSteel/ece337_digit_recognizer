// $Id: $
// File name:   pts_shift_register.sv
// Created:     4/4/2018
// Author:      Chan Weng Yan
// Lab Section: 337-08
// Version:     1.0  Initial Design Entry
// Description: Parallel-to-serial shift register
